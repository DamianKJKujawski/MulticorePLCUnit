module PERIPHERALS
(
	input 							CLK,

	//IO:
	input wire 					BITPERIPHERALS_READ,
	input wire 					BITPERIPHERALS_WRITE,
	
	input	wire	[15:0] 	INPUTS,
	output wire	[15:0] 	OUTPUTS,
	
	// ------  Bit memory ------
	input wire					PERIPHERALS_BIT_EN,
	input	wire					PERIPHERALS_BIT_WE,
	
	input wire  [15:0]  PERIPHERALS_BIT_InADDR,
	output wire  			  PERIPHERALS_BIT_InDATA,
	
	input wire  [15:0] 	PERIPHERALS_BIT_OutADDR,
	input wire 					PERIPHERALS_BIT_OutDATA,
	
	
	// ------ Word memory ------
	input wire					PERIPHERALS_EN,
	input	wire					PERIPHERALS_WE,
	
	input wire  [15:0] 	PERIPHERALS_ADDR,
	inout wire  [ 7:0]  PERIPHERALS_DATA
);


WORD_PERIPHERALS _WORD_PERIPHERALS
(
	.CLK(CLK),
	
	.WORDPERIPHERALS_EN(PERIPHERALS_EN),
	.WORDPERIPHERALS_WE(PERIPHERALS_WE),

	.WORDPERIPHERALS_ADDR(PERIPHERALS_ADDR),
	.WORDPERIPHERALS_DATA(PERIPHERALS_DATA)
);



BIT_PERIPHERALS _BIT_PERIPHERALS
(
	.CLK(CLK),
	
	//CONTROL:
	.BITPERIPHERALS_EN(PERIPHERALS_BIT_EN),

	.BITPERIPHERALS_READ(BITPERIPHERALS_READ),
	.BITPERIPHERALS_WRITE(BITPERIPHERALS_WRITE),
	
	//In:
  .BITPERIPHERALS_OUTPUT(OUTPUTS),
	.BITPERIPHERALS_OutADDR(PERIPHERALS_BIT_OutADDR),
	.BITPERIPHERALS_OutDATA(PERIPHERALS_BIT_OutDATA),

	//Out:
	.BITPERIPHERALS_WE(PERIPHERALS_WE),
	.BITPERIPHERALS_INPUT(INPUTS),
	.BITPERIPHERALS_InADDR(PERIPHERALS_BIT_InADDR),
	.BITPERIPHERALS_InDATA(PERIPHERALS_BIT_InDATA)
);


endmodule 