module BIT_PERIPHERALS
(
	input wire 		    	CLK,
	
	//CONTROL:
	input wire 			 		BITPERIPHERALS_EN,
	
	input wire 					BITPERIPHERALS_READ,
	input wire 					BITPERIPHERALS_WRITE,
	
	//In:
  output wire [15:0] 	BITPERIPHERALS_OUTPUT,
	input wire  [15:0] 	BITPERIPHERALS_OutADDR,
	input wire 		 			BITPERIPHERALS_OutDATA,

	//Out:
	input wire 		    	BITPERIPHERALS_WE,
	input wire  [15:0] 	BITPERIPHERALS_INPUT,
	input wire  [15:0] 	BITPERIPHERALS_InADDR,
	output wire 			 	BITPERIPHERALS_InDATA

);

INPUT_REGISTERS _INPUT_REGISTERS
(
	.CLK(CLK),
	.INPUTREGISTERS_EN(BITPERIPHERALS_EN && !BITPERIPHERALS_OutADDR[4]),
	
	.INPUTREGISTERS_LoadInput(BITPERIPHERALS_READ),
	.INPUTREGISTERS_INPUT(BITPERIPHERALS_INPUT),
	
	.INPUTREGISTERS_InADDR(BITPERIPHERALS_InADDR[3:0]),
	.INPUTREGISTERS_InDATA(BITPERIPHERALS_InDATA)
);

OUTPUT_REGISTERS _OUTPUT_REGISTERS
(
	.CLK(CLK),
	.OUTPUTREGISTERS_WE(BITPERIPHERALS_WE),
	.OUTPUTREGISTERS_EN(BITPERIPHERALS_EN && BITPERIPHERALS_InADDR[4]),
	
	.OUTPUTREGISTERS_LoadOutput(BITPERIPHERALS_WRITE),
	.OUTPUTREGISTERS_OUTPUT(BITPERIPHERALS_OUTPUT),
	
	.OUTPUTREGISTERS_OutADDR(BITPERIPHERALS_OutADDR[3:0]),
	.OUTPUTREGISTERS_OutDATA(BITPERIPHERALS_OutDATA),
	
	.OUTPUTREGISTERS_ReadOutADDR(BITPERIPHERALS_InADDR[3:0]),
	.OUTPUTREGISTERS_ReadOutDATA(BITPERIPHERALS_InDATA)
);

endmodule 