module BITCORE_ARBITER
(
	input wire			 		CLK,
	//Carry in:
	input wire			 		BITCOREARBITER_WE_Prev,
	input wire			 		BITCOREARBITER_RR_Prev,
	//Write
	input wire			 		BITCOREARBITER_WE,
	input wire			 		BITCOREARBITER_RR,
	
	output wire 			  BITCOREARBITER_RAM_WE,
	//CORE:
	input wire					BITCOREARBITER_CORE_WriteDATA,
	output wire				 	BITCOREARBITER_CORE_ReadDATA,
	input wire	[15:0] 	BITCOREARBITER_CORE_ADDR,
	// -------------------- RAM --------------------
	output wire			  	BITCOREARBITER_RAM_WriteDATA,
	output wire	[15:0] 	BITCOREARBITER_RAM_WriteADDR,
	
	input wire			  	BITCOREARBITER_RAM_ReadDATA,
	output wire	[15:0] 	BITCOREARBITER_RAM_ReadADDR,
	//Ack:
	output wire			 		BITCOREARBITER_ACK,

	// ------------------ Carry Out ----------------
	output wire			 		BITCOREARBITER_WE_CarryOut,
	output wire			 		BITCOREARBITER_RR_CarryOut
);

wire 	 _WRITE_ARBITER_ACK;
wire 	 _READ_ARBITER_ACK;

assign BITCOREARBITER_ACK = _WRITE_ARBITER_ACK || _READ_ARBITER_ACK;

BITWRITE_ARBITER _BITWRITE_ARBITER
(
	.CLK(CLK),
	//Carry in:
	.WRITEARBITER_WE_PREV(BITCOREARBITER_WE_Prev),
	//Driver data:
	.WRITEARBITER_WE(BITCOREARBITER_WE),
	.WRITEARBITER_RAM_WE(BITCOREARBITER_RAM_WE),
	//Data:
	.WRITEARBITER_CORE_WriteDATA(BITCOREARBITER_CORE_WriteDATA),
	.WRITEARBITER_CORE_WriteADDR(BITCOREARBITER_CORE_ADDR),
	
	.WRITEARBITER_RAM_WriteDATA(BITCOREARBITER_RAM_WriteDATA),
	.WRITEARBITER_RAM_WriteADDR(BITCOREARBITER_RAM_WriteADDR),
	//Ack:
	.WRITEARBITER_ACK(_WRITE_ARBITER_ACK),
	//Carry out:
	.WRITEARBITER_CARRY_OUT(BITCOREARBITER_WE_CarryOut)
);
	
BITREAD_ARBITER _BITREAD_ARBITER
(
	.CLK(CLK),
	//Carry in:
	.READARBITER_RR_PREV(BITCOREARBITER_RR_Prev),
	//Driver data:
	.READARBITER_READ_REQUEST(BITCOREARBITER_RR),
	//DATA:
	.READARBITER_CORE_ReadDATA(BITCOREARBITER_CORE_ReadDATA),
	.READARBITER_CORE_ReadADDR(BITCOREARBITER_CORE_ADDR),

	.READARBITER_RAM_ReadDATA(BITCOREARBITER_RAM_ReadDATA),
	.READARBITER_RAM_ReadADDR(BITCOREARBITER_RAM_ReadADDR),
	//Ack:
	.READARBITER_ACK(_READ_ARBITER_ACK),
	//Carry out:
	.READARBITER_CARRY_OUT(BITCOREARBITER_RR_CarryOut)
);



endmodule 