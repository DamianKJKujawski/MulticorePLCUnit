module WORDCORE_ARBITER
(
	input wire			 		CLK,
	
	// ------  Carry In ------
	input wire			 		WORDCOREARBITER_Prev,

	// ------ CORE DATA ------
	input wire			 		WORDCOREARBITER_WE,
	input wire			 		WORDCOREARBITER_RR,
	
	inout wire	[7:0]  	WORDCOREARBITER_CORE_DATA,
	input wire	[15:0] 	WORDCOREARBITER_CORE_ADDR,
	
	// --------  RAM ---------
	inout wire	[7:0]  	WORDCOREARBITER_RAM_DATA,
	output wire	[15:0] 	WORDCOREARBITER_RAM_ADDR,
	
	output wire 			  WORDCOREARBITER_RAM_WE,
	
	//Ack:
	output wire			 		WORDCOREARBITER_ACK,
	
	// ------ Carry Out ------
	output wire			 		WORDCOREARBITER_CarryOut
);

wire _WRITE_ARBITER_ACK;
wire _READ_ARBITER_ACK;
wire _WORDCOREARBITER_WE_CarryOut;
wire _WORDCOREARBITER_RR_CarryOut;

assign WORDCOREARBITER_ACK = _WRITE_ARBITER_ACK || _READ_ARBITER_ACK;
assign WORDCOREARBITER_CarryOut = _WORDCOREARBITER_WE_CarryOut || _WORDCOREARBITER_RR_CarryOut;


WRITE_ARBITER _WRITE_ARBITER
(
	.CLK(CLK),
	//Carry in:
	.WRITEARBITER_WE_PREV(WORDCOREARBITER_Prev),
	//Driver data:
	.WRITEARBITER_WE(WORDCOREARBITER_WE),
	.WRITEARBITER_RAM_WE(WORDCOREARBITER_RAM_WE),
	//Data:
	.WRITEARBITER_CORE_WriteDATA(WORDCOREARBITER_CORE_DATA),
	.WRITEARBITER_CORE_WriteADDR(WORDCOREARBITER_CORE_ADDR),
	
	.WRITEARBITER_RAM_WriteDATA(WORDCOREARBITER_RAM_DATA),
	.WRITEARBITER_RAM_WriteADDR(WORDCOREARBITER_RAM_ADDR),
	//Ack:
	.WRITEARBITER_ACK(_WRITE_ARBITER_ACK),
	//Carry out:
	.WRITEARBITER_CARRY_OUT(_WORDCOREARBITER_WE_CarryOut)
);
	
READ_ARBITER _READ_ARBITER
(
	.CLK(CLK),
	//Carry in:
	.READARBITER_RR_PREV(WORDCOREARBITER_Prev),
	//Driver data:
	.READARBITER_READ_REQUEST(WORDCOREARBITER_RR),
	//DATA:
	.READARBITER_CORE_ReadDATA(WORDCOREARBITER_CORE_DATA),
	.READARBITER_CORE_ReadADDR(WORDCOREARBITER_CORE_ADDR),

	.READARBITER_RAM_ReadDATA(WORDCOREARBITER_RAM_DATA),
	.READARBITER_RAM_ReadADDR(WORDCOREARBITER_RAM_ADDR),
	//Ack:
	.READARBITER_ACK(_READ_ARBITER_ACK),
	//Carry out:
	.READARBITER_CARRY_OUT(_WORDCOREARBITER_RR_CarryOut)
);

endmodule 